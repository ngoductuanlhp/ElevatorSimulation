module one_4_mux_1(in0,in1,in2,in3,select,out);
input in1,in2,in3,in0;
input select;

output reg out;

always@*
case(select)
2'b00:out=in0;
2'b01:out=in1;
2'b10:out=in2;
2'b11:out=in3;
endcase
endmodule
